//Logic Gates code in verilog
module logic_gates(input i,j; output 
